----------------------------------------------------------------------------------

----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ctrl_unit is
end ctrl_unit;

architecture rtl of ctrl_unit is

begin


end rtl;

